
module InstructionDecoder (
	instruction, 

    	
);

//Inputs
input [31:0] instruction; 


//Outputs
output reg [1:0] firstLevelDecode; 
output arithmeticToSpec; 
output reg [3:0] secondLevelDecode; 
output reg [2:0] aluOC; 
output reg []



endmodule